library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.psc_pkg.all; 



entity fofb_top is
  generic (
    SIM_MODE     : integer := 0
  );
  port (
    clk          : in  std_logic;
    reset        : in  std_logic;   
    gtrefclk_p   : in  std_logic;
    gtrefclk_n   : in  std_logic;
    rxp          : in  std_logic_vector(1 downto 0);
    rxn          : in  std_logic_vector(1 downto 0);
    txp          : out std_logic_vector(1 downto 0);
    txn          : out std_logic_vector(1 downto 0);
    fofb_params  : in t_fofb_params; 
	fofb_data    : out t_fofb_data
  );
end entity fofb_top;

architecture behv of fofb_top is

  signal shift_q               : std_logic_vector(8 downto 0);
  signal fofb_clk              : std_logic;
  signal fofb_rxd              : std_logic_vector(7 downto 0);
  signal fofb_rx_dv            : std_logic;
  signal fofb_rxd_dly          : std_logic_vector(7 downto 0);
  signal fofb_rx_dv_dly        : std_logic;  
  signal fofb_txd              : std_logic_vector(7 downto 0);
  signal fofb_tx_en            : std_logic;
  
  signal fofb_packet           : std_logic;
  signal udp_rx_done           : std_logic;
  


  attribute mark_debug : string;  
  attribute mark_debug of fofb_params: signal is "true";



begin

fofb_txd <= fofb_rxd;
fofb_tx_en <= fofb_rx_dv;

--phy instantiations
fofb_phy : entity work.fofb_phy
  generic map (
    SIM_MODE => SIM_MODE  
  )
  port map (
    clk => clk,
    reset => reset,
    gtrefclk_p => gtrefclk_p,
    gtrefclk_n => gtrefclk_n,
    rxp => rxp,
    rxn => rxn,
    txp => txp,
    txn => txn,
    fofb_clk => fofb_clk,
    fofb_rxd => fofb_rxd,
    fofb_rx_dv => fofb_rx_dv,
    fofb_txd => fofb_rxd_dly,
    fofb_tx_en => fofb_rx_dv_dly
);


--FOFB receive fsm 
fofb_rcv : entity work.udp_rx
  port map (  
    fofb_clk => fofb_clk,         
    reset => reset,	
    fofb_params => fofb_params,
    fofb_data => fofb_data,
    rx_data_in => fofb_rxd, 
    rx_dv => fofb_rx_dv, 
    fofb_packet => fofb_packet,                                  	                         
    rx_done => udp_rx_done
);
	 

dly_packet: shift_ram
  port map (
    clk => fofb_clk,
    d => fofb_rx_dv & fofb_rxd,
    q => shift_q
);

fofb_rx_dv_dly <= shift_q(8);
fofb_rxd_dly <= shift_q(7 downto 0);
  







end architecture behv;
